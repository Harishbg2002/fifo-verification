$display("WRITE: %0h", din);
