// Driver class
class driver;

  task run;
  endtask
endclass
