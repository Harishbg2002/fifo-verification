"// drive wr_en"  
