hjbchbvjbdjvbdj
jbvjdbvjwvbew
vjnwkjvwkjvb