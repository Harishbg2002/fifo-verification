"// check data "  
