if (wr_en && !full) begin
  fifo.push(din);
end
