jghgkgdkjghjhg