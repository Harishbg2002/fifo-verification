hello world nvkjnvkjfnvknv 123