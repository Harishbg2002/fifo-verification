hjbchbvjbdjvbdj
jbvjdbvjwvbew
vjnwkjvwkjvb kjnkjbb