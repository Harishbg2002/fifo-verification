"// This is monitor"  
