// test code for under_flow