"// This is scoreboard"  
