Command: git pull
○ Fetches and automatically merges changes from the remote branch into your
current branch. Use this to keep your branch up-to-date with others' work.
> git pull origin main
