hello world nvkjnvkjfnvknv 