hello world nvkjnvkjfnvknv