<<<<<<< HEAD
<<<<<<< HEAD
"// drive wr_en"  
=======
// Driver class
class driver;

  task run;
  endtask
endclass
>>>>>>> 72c8ae165bb4107438102f54f7c4a4ffbf2b7f57
=======
Command: git pull
○ Fetches and automatically merges changes from the remote branch into your
current branch. Use this to keep your branch up-to-date with others' work.
> git pull origin main
>>>>>>> 807ef19e586eef052f5abcb6c16dcc51f8c24d83
