<<<<<<< HEAD
"// drive wr_en"  
=======
// Driver class
class driver;

  task run;
  endtask
endclass
>>>>>>> 72c8ae165bb4107438102f54f7c4a4ffbf2b7f57
