jghgkgdkjghjhg
hjbchbvjbdjvbdj
jbvjdbvjwvbew
vjnwkjvwkjvb kjnkjbb
